// simple and in Verilog
module simple_and(input A,B, output O);  
 assign O = A && B; 
endmodule  